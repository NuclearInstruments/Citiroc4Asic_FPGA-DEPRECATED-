--This example file is for demonstration purpose only. Users must not use this keyfile to encrypt their sources. 
--It is strongly recommonded that users create their own key file to use for encrypting their sources. 
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
JwXK2b+hpdQKCG/aofkd3lHFK74YnjI5wLLsN5G2BIqIQ0raCicqceEzXCRDwNtVHaJ6UD66WZu8
w/O8XimFFXHYUeK9Yg8oOkAfD7H0RBMathr7RLH/lQfhyLFaa1N0b5cfLCSsJdHRRqIhCGjA30AV
gYag+RjfxN1ehV7wbQOGXhoHaUcpY5ttx3CQkIkXpHNyG5NzAYqxGubXttoTsRElEqJINIKRGJ5O
XKh6LQ2KzQWhcg8a5evGxd7qXrfDBF8acf+3ndqpHux+LE5H7SVd5V3D85LHfS2gXU8msaLFqFWD
X/WpOLQi9yJ+0MTeH3bF9v8bpcKExaeJec5UPg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="1fRWPTCdWTHe3Jj4jaalGamNhHykUs2j8O1aTbwiKK0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 27184)
`protect data_block
MsuhZVg/FqeDSXiddbv816yMwJsgMYnqsXGyTyUudJm7aatlGsWEeqFl4F4LML8DLgkRefuagqww
vndf+v1lP6GGrogVytwnCCkknZu4kHphAuwpbk+RJrX52eflKL2kRIfGUo7THrYKUpFnEfo2YEqA
/U6Wh+LvNFNYERvDJjovmqh79dS54dawL4a9lrTzCLliB/OilDDh/NrezXI6+4aU1HELYVAsl2Zq
vfjNPllUiEvIBrboWhqkCeCOU6S6jiV6uVnl3+TSBGXP0Y1jU7+Ksk1mrV0kbqs4fF9MvhTmaiRK
xpC5CRW3+0dA6VXKPIRL2IQ786SmgJMmQo1MVlC9WWAESrccY4TXA3A++ls1TyaW6Y9609xgqSXx
3u+//B7+4/88lp0RPbIFZ7i6MVxsch4w2QY8o9aRH+9qPYcSp5QE/3uClbfOC7h3E4erT2JP2/B2
TArAVTKRUBp6eQ1705OBMBR9n5aqhxE4BNh90LQOL1puS5hpsEndntsAiT7VqDZmvlb0UFM08pa+
e2Jy+Uo83kI4LAM2o9mx4DOKBueoWx3nuWfKt8cKI4CL4poLOUe8M8fProKyZKgKlf7ra/Ess0Jf
WUWvI5vLlYoEkd62WfJatVk7MCjZM+fcklcBuujPVPDqg+O01HOdLwCU219X6VEq82ZjvwCyZFA3
PP3xN8SRsabYtnKT+0yXWNWzM/tNy9Tuaj0ABUVJC7i8+WHFv82W54YDbcDPwUn5PdIthmVjq+na
i9jxC2Up6OW6l7AlY9USkPVCekHqseZCtlH1HBwamQrlWZqwz0YHJG4ok7rXvzrjvCDWDgfZhU93
UqryS+D5ehzCTVPjMrmTCgA68cWjNBdkcz9gT8LDcpU7LMcZT7nfYf2KPrWXRDisiD84DQDyOowL
aOpfLKpjbBiqALawn4+YRK6rHb2bz9JVNoRKlmzq/GGY1dYviffS89cm0CaLmeJMAKRK9O5tmPcW
ZJhvKcq3Tpq4MrvFLLrmt/KR/ST4pGT/4p1CX/JwPfuLR6YwWkFSeqKChumW18IwcEFpeFjQVLoB
UfMvKc5AiVeFmI8EcffJUJ/n7uZiGK9arIHQZjj/6uHW2N3GfkEgm0muIm6l6l50wFGZuluSTA9Y
zLT5hp3a07O/fTekOf32E26H/lEMwPVDnNHPDhPrzdAR+ozJJnhYllTrhjfm0v0yvp7IkuuQiIy5
3MgYdDKghrILWQ6ovr0dIm93RawsLXhkpcYAF4Oa/6pilyv9XPE4MJT5zYmzV86FLyXmnHe691Jj
utHkmvpzXu0DJDP8DUIKCE9CE1/5nFmMG4hIFZTi1h0Fj6gsQ7I2gYFKy9EpXqzNuQ6DHkh7dX4l
kw+w1RpTPt7oVJhtzPSH0L2Oo6zVN7Q5qWh8IY2B2/Ew93IPOsTg5XJNh48ZP95goEMeii9mB8aS
lg9bYj5sCv+OGC0HMOgWju1V2Jfy4fWWmjj558o8bCyw3c5qpVyKbG1sC/sND+xLI8F9WYgAFlij
NgO7+N6kTeuH7f6OkY9Y+ff02PRe6ZtMIFMFP5vcIAZO+sIilWyrK479Vy720tqXumxjOnTsNgWW
y9dWs1gMC19MtRi63kujzEUFm5tihIc1ng/GN9bM2+EacAnag9mVSiqh+70czRXW3HHaR00fQZM2
Dpu4Y+hFIxo1B0NVpeyghlBUmcG5AQ315W5Pnp6dmQbN38T838dz9VIr79M1jzY573Nv+0EaeGTO
RKm6/jqqyVs8htW/ljgd0Cvx+etPbBP13t1bwJW0bPpK8X6r0aeL5L00k982TYNFMn3N0B+om18l
r7Yz9LG0zBOenp1go9xwLo/YEam2u086Awdvd9z5EuuEezRZWTGbTe23Xp+53X5loU/VtCmSj7Ap
iR7b5Cn0WSDLgcdkpDdTmWp5bQKuYopNeew58FZFz2csUf5h/7tujrxOb2cvSjC6p1Gq0MZd9RmN
U9K3NJFsaJdpwbZzPcWehabfEqLvMrP5RRs9kr2QLLNG1jdvgAMiq4NFQ5AqLUbCSZCmoYRc2JHR
dRu7Azwl1gY/7nBpd5sEDlvd6z3/yEc3gf3lNpg7vCoJj2ekU6Ykh2ctCUm8phIlwMOtN76R6OEb
tfW1PGfdIGlhKNd6Wt5nFA9vEFbDICmbX8O6LxO90qLwKPtO5hHGD/iwBd34d+Vfgzuj+gZCi57A
Hvj94Ql5rD1GEXoMnzrKNAHBwp2QcgXm6VFIn51GqeZvImRvYYqeLQFg+HvFjWVWZjs8fXzZ+aZO
xvRbbcD1JOHSwD5zlZVI6r9G7RG0gAqJEMA2FmTZzuQaAEVXThssWxM+gqwBfW3bisTeoQ7/5FhN
XyomRf3rPWQF9UWn3P63oguJGDHLsacKfGB5zlussDB8NtpXxskXgQQWDW5OFB325QMF930n6/Uc
G62W5eZDAvJHml3ntIYsnwlmMLidG0DInKGTx8SOj7whiB2PVIiAokKmr27hHxwnJou9HTp6+N5d
RLnA5EDXwodaEZFfpHJa2Z5Lx1XtYCXojlHUcchz6is36AyQZXPJ6RtyrZl+p/MWH03p/u8xLJDi
vEHvGv/m1hsJfa1pfH4c26hRiWysSyIacI1AmEl2d82VXPUXasN8C2tbAIk5FTRyOhk0WEVQVcXG
9j9hdEiwzpnpBZD9teO36+K+/pHs1VMjVRNIB/RdgCk/OFwUpX0UrkO4do5mqoiqXiWMxqK67pAb
wx6oCSpTm3oM9HbJbYtdGaOMkl4lqpwYZAGKnMqKGttzYpXfr45X3I8QKWblY7XMWxpp8nCf612I
rqqEwR9O0eHxXOyjoo8DgpJNe00qXclNSDaE6X2LmoPiPKzSG2t6jq+VDg2lrPkWn07u9udBXV10
AYJ9wHz/OvpIg1o/zPImLZuaLcRZqr65MhJRhma5mw1pQz1nHLdJA77hXYJBfPmtobAX7IFGSwjX
gNkvcaWlYUTNdH8NYtjUC9ZJZBs4TTh9dMqSmTUizXNLdweIwueWi7IqQRG8ecqOQRSuNVq+TUTz
V/LPrZ3gNNhOXTljx3bZkovQKbN7i4hcU9kE1D2jBndm6DDErF4Pf39tlWyovsvtjKRPOed90HNg
57X+37BbcPxs0syvX52yhIsy06cFh8mzxufig71jwK8yDM3Vi9PEUwvbiHQzTO1SR5jHplUdh/tY
q91SYOzT28KQSQ8AKAuBPaLLA4FNk/fqfafBnlxVqYpIBTCM7Ebzvj6dy6dSAhpbWjqx4Zwma2/q
guRQpqSYhDWi2tMtIN29w9oBDRz/5ppOP+pmqGEaFSoV5CtKRi30D0TUtKIIXrCQjX+zJJi+7wl2
h5me2I7UOdorYP0r4Ob8TROVuwB+/3p+bncJj5SmkV2/CiXtP2pBnY9NFkHX6l1/MvfPivMecTvP
9WenixphJwlGhpdHSxixddoLCLZSU7gKqBncxy2Mnyg74vrdtLf7Ae+3IleciqiBXCOIeuNlptKR
Mx6W1cwaMK9c2H3pbuo80R+Cr8QVJ8SMRuqDXsq52rau2xGUC8NEBfzmHwS2CVWZ//54bGbVlo8S
8V+1TiphHpG/8WnBjVzwnU0ITCL+tgLViSdEOMzotB1fBLQvn8L2g9lpnaVzr9WnJ3vCvrwIXCd8
Z6JSXRBla3I81gjqOgksdv15geICRpG57cFMBq5R73u6wi/VLwd4v27xG1068Bz0xgDd+5jOTOlM
hvx6IGpRlMzIMRJLWcccnt2SBWBY5ZFBAqVwkM4DExzAntQ6PaLCc736Ub46qCd8v3rtNyM4IBRK
36iQCJHfXjsd2rdEYj9PysQtgpfoO+G4GnNeeQMZ5A1uUV27ArIUaOg7UGPRxLVn9En8bPuIgEop
e11lI0iNvD6iksBgx/EGaPRYFMe98M54ZK52PQjUPjJyc89lV509nYV1jLworfgFYij3T8pk/QEH
EQi+A+3wrhXma4RVyzpi77Nnp118pzdwTNSXFCQ2MZygyGIniA6EKK1ooxNn6BVevdxI1LqdYJ83
FQRdsbgQfd8RPk63WcM9n6T4yCovgQuztEyzyIirZf1mR3GCbV7IzpvoRyvPwhrk33fSi4ItW1+D
eKClSAASzgKKc0Zywrh3NPI148y1H0hN6wA5qVvOw/c8d1s3EP+pS/Pb6urj8FyXbWEJ72uiq1Ax
oWvJccSPzZgqzWtpzq9ZMt4Kd7I1csUWqRf20EoC2FZfsfHPP9CGJK9ZF6IczsEfH9uGntEh9Dfy
wu5ZYiuJ7atDuOKecyk7nN1QSjF28sLDDHqXssQPhY9eGkYUt5WYDTma3GK1pKGSpc5ghPDUA0f3
PWalwAhEcN3NuEIRRmS0giW1eczrBDhU0yGfdCtE+GXHFN6rpDUQn/hD+DSo2F7R3in2qRUjIepi
BOvL+s3H/geBlTs6juyeQWUhFefG0if725I2UWjYauwWx9y2QO7GSbA2hBEqFhJbqkCdYb12BJlx
rdWpQ4T3PYOY2lZF083TGr001KRgRuZsvpEolNPTwSO12KbIsVkgZ/YNFESBCgv+Hxk0vmF/pSWD
sBBC+zRDZ7OFz8NQymNL9iWRPH+bsPwz1FdAr50prsmQUzhvyRaVRRa1pnETb5waD0UvwLFwYll+
IGudttVqOl8mKSReRdl7Kiq6K81Eq61GTlwCYadCm5OSXXnWg+6PdMjkGbssOnH15Vj4tJU934gj
dvZrWzrUwJ50bXiwpnHHFAuDACTxrUZrY6t0MIRMipqzdWxCG6nLOsMb1G8dFGaS5Rvc31tWIgKE
HeUWZPrS09MZp5zfQpTvSdgh6cBsK/Lci9o5oBNcCQs3wg3zVKQpW6AtiSFi44NmPwu+rxRLGpuw
s3a4Cp9pQGejGI3EhhRpNlKAZtwCc5RcMzisG1yxngxpef6GWabBN7yyzmM6QRwslr//X7PWMKdn
YkFcXfXxqtC1tlD8/mYNfcDauCRPDgDjFmbXv6QZDzck7j/ixHAVfR7DVDmplfYfvGYR0hNzLTD9
vMDJaw9vmrER2B7pwzvb6LTAdNYxNk31gSSOW9QCP9LzRg4jtFRWVj6mXnGmNME1vFQfYwRvkdaB
nOzsE1WfsmONmcFICbjywjkRw4eHmSjGPyQokkgmmce4bIDS/aeD6TuifMSWhZNsYfvaA3ipa3Hs
AK4XQIR05tmjLG9MulAtJDdCppi+Xc4qgbh8YlCiNKyhicEkSy+PJZ/o5cLfbKHsNeEMuXdSCtoW
mJSnqEXCe77vzU9cGVdkp/RJiVs6n3y5mny3Axc9EG/7xn4oq9l2oFNNTG4Kaz9DSj7WNEAy2Iw0
iL3rLvklMtkMtcR8CzfpwztmphkXiPEGmrDGmNeKke7ov8RmZa00WAiZZNO91Uo6imrfXv6Ntl7Q
1CMsEkNCjmDh9O1uRUUDFjOnlPtq5kM+Yn3BtmzzKWQv4Ou451repgSp6FHOOnRmWA7C6jdby5nV
v9zIHSh/G8cXXcmcNZH9jsQ74yNtBwdaxAKtGVUjv/7GL7wtNYu/Vo9AiAPeL9BrIQdDAwZDcaVr
9oyF6qfr5y8R4AG8P3Bko+FrpH4JzLHtsyBGxR5b0esEildw/69rfM6wMsSV6iIsO6Z4cmat57Ag
i+WrCTcAtAEUpQtt+/DUqIrjGheqmrx0m3qBTyRU3aoBRF4EB3A7dCR3xd0N3XLET1k7jmTzVM82
JbmnRONjCoasvcFqFJFPg+eysTWmBwDIOESoEVQsvMiK3kIYf54bgfZIS9osfyRt5vTiqbt5QumS
DL7vexh+snvqwCf11zDEMIQSCl26PZxieh6TWHJHPhrqdDkVd6rGPwWc3SRBD290ZwHLFh68Ncz0
ab3I4ViKK/vlbrqR8SNa8EV3kQCDvvaQqf13lGDKEsmlz5r4dspdngT4nNZnMaWYouTpkOLv6r2J
gC+TwqtV7PaDMnSlApdPqS1DZWSKwXz9m/3nEqT6if3DD57MfYk3KyXdw/NOBkmQpZz/09UOmlmf
Qpmvwm8Cj2VHgjS6SkOcpaWGBN66SIWm0a7gz6fm64LPgUXdkfMfTP4wooUAaQ3W/mDWBD7tG8Av
+vCweFtbjhMQ+LQMd7ai1A6gCCedqyJrWmcF2uwCstDdxE38xk6nUP2KRdLqrLwCk6BddYMZoXUU
zRzZLxiSfO3PsuwYlo2QG+JCve+3f0ruk8md4GIDFR4ArXB4nd6Jlj7ZRMSfdUzlj1oKO7FRM4o1
WUaqz8iKuJrnUoWVxH5pNvZJ4JSR4dvbpWhXDoQy6CikkzTLZYxD2dVpeA5Ct9TkL2J2NVyZqCNa
52O6RfEx80yenGsXTFEZSeoMJRBQrlVhCLQ6UFHub3W+QuTG/cXhAM060RWAdVT6okXidX1T59rf
FVDb/zdQQRR9El4qV32Otckd/fYeDc9lFXCCjz/8DnjYFo/i2b8sb0YQcPHAAX3AKyLG/qPXVl7t
Fz+kJaMt/mvYYQzXFRtZ1SBuNhg1riaYw5MFw1Ebmr5gAEZTEw2bmNY5ahbuXeVb9dUJjIxzwYjn
gcVMWQsQ+/2M6GZ60B0LSaJhJBeA4bKkM9b/cdzpwBfweHz0GWNdj8BkTV007hBPtTRagr9GJGtL
h/wfTNr8xutoY68kd/6lI59UZvBXadPiXFyxed0lsEOk7h7HX2L3AfjF502VyK8q+otrU5peODTY
z5oAhC+iPeusFVi3woZak+B4tO4KevxxCDDmLpilaqVEtU9nG+4ibVl+9dwoWiR4Q1o0m2pQ8qOV
VH76BWN7JdGknCR8zXDVwvNVepwsn4yGYkUer3f3aDu7oB6X4mKhJzO2UmclVRUt6QF/AgIuygqc
ijTSrgAkWu17NX4VSmhSiVh7eufgN/yqoTPkUMwsty4vnuyBvE/OibFRvzY5NecKsf2A9DNzWrwP
8P5WhfzBe2yOaAo8Z+GjMLuziUSVWLt1Pd96WCfHSghoHLlHywzAS2O6flqh5m8xnK0frsgfKm0F
H5k8Mu+hd90KMjy0aYjItg3HCNkpvPais/+2oGicWzrwgardk+zLad4HRGf97G342MFbbl/7ia0C
2SL33/2VDiTMdrnJFxLTdmCMVh25ywYoS6ME02k2yLF7kkp2EQOml7bMOPF0M1YfgcsBci8WA0A8
EPI5HWJXXMe48YZDnyXE/cKzd2iUwmzXQnJqxIig9zbzgQeyVOvjElcbdM8n3q0tJ5DkwP75xeD+
hPpWmAcKyertpyRI4exaKfKHxrEltprKIBD8e7aJ3JjwyHRA9TL+95bz73G2RtqaSX6KQXAhVMPO
eycCExPYFa0YRX3whZbIeLpFc4va+YnVgqyM9cNhDbTdpkRHBu15RDSddBm89UOU3ClX5OJUx38A
dvFRrNG9XXHLkd7szOZvR8FgvVeB5nIAz7pZGGtnTZO9/NkuQpEHCII0x/YFidiFY/8dTO/QowND
mrkIv+pbrLrERJd2D6r/MezY3vpStRVQbPvQHKOhFHg0B3N/3NnOP5da/HI8FixnIlruw+/t0Ban
eqj+edJKtiyvp8Y8KpcPzbWDH6svFr7RbiVUHP4BxzapSvcP7q3z2poFnP9ikE0XqDBuQntqm8ka
hS2L/QDS87lS3a6mBDbPGVMdMrYtcCxJmTOfXNz6xhHuAgreKDBTE+BdrrZ2m2SDMvNR5X2w3ln/
KFgZ32YjPL8AClNCAp3iEDMGg5RwVQNazw3+svzcKDNYm+jIlnRmYHSRLk/tGaMHwuw59hxk4m8Y
+aoEr3a6FX5vW40Tu0j8gyX/rFd1sgrWgGD2jMT/dJFWdp9Y2NGrIZA6iNWx7I90SpbasDouw2tU
PX+IQNFqdYyfVmd0YWJ7fQG6iBQg/IxtgdFrNM6t+b4uYPgz5R3mVgOqL9sLUj8BO8EuATsttKQe
mdEnnWiXVYrfV15gQUi9V+D2M5ovqA+sj2Z3YFzE8Vd0dIygTn6DK0l5nnFhdpjL5meMkUHqLTx6
bwVHETCHapgRkEcBTwGM3lGN2ZwYDGkadD9GItQff6wU+WvgejcFIOSB9kY7OOC10zuRdGH5GGZW
h1zBE/vIH0Cxbr6QAs6MDRzieyjITSKaDgUpM+GQcUhD4j7HoO/BwC3KSAdxF1b6CEocFle8tcqH
z2tNu2/U3zweLnkJgn6CMAkUWervmvtQ1yABLqnhHB8VfBFWnp0ToZxXv65Uk5QXIYK8WxaymZP7
u1oKePLoPlER6pxcnfKS+oR3z48XqFnSvS+vHrKqqR8xZhuhpqUtptj1Ha6JZRe3Giimai5Wjtdf
y1zb8Lu1/lEllrcJDEI3TaBhgOwS5J3aRpTWICRoeMa9LHZZHOmOkJRguek2graC+jKPmLO3ZmbY
RgayLNrjXYbf5MZr/pkMhNvZWjViS9wu/pvVYBCHYem/qIOub//jM+NqOs/87piS1F0PGRuNkqNK
s1sw05Dke74xztujp8bMsl6MiXfKeYK3yJXU+eb7iwavsVFlWMRvLE1ddX2I7+LJ4P2eI/ZMVjQy
Cwso8smP840G9JyZXIiW44HdcyyN6IL3yMDhDrSE66scdGgh2mOVmwk4opfsQaKMXTec3cqdimNv
bZ3W3/w2cpteeE/Xe4o7ztizRJwCfOD4ilAQsI9WLP997aR+hCokmjn7h0BvVfFZh3NKubDmwr8j
ZZiJrTHXF/YR0KtvAUbpHZi/BAoWqr0u86ouXNRxvbhRra9Moem+wAyPDr/ls6FfuIFE24BDNZQQ
M2xHk0849Uol7aCuuhwB1KbW/ZtlLZhCq6UllbwFvUz69k8cJM+S2olN5nxqa5fVbzOrPsWjPUVJ
G+lTfR2lhl2d8zx6ywqcy8bOd3jhetXBHJY6Jd7KxaRbUgfxDCuy798LF1e3cj4Xi1OvTUBhXfXy
c6RMjlXB0viFzFEnl5JN1m6AdYMZ1JV5ObUjXwIEnAUMnrVKdAO1nzNGeuO39CvgQk5veH5h/p+6
LU0ce4NZ0FASLu6T9Bf0X0+9UNpjv+y8zYIseJfJGJ/3HQc+vi3RA97dLMPnGXUB3PXwMuvngDgK
jYu+xm41MT89yH+vN7kxWjczk0hssg7cte++jK+KD/VCIQRtDAagtJgwNXx4mgHYeeUq+J/jt4V0
X4FiBbADpZDzVplCvEdj3/oXLFX3cIN+VqL6nK8DGDMIXs3xZIIszIkTapZY13XA+9KSN41gx8Yk
poolWrjJzaX6vfEcwwemtDFDIa6/z26QqatLZIp/wkyQP7d5fWoVWPt3Tg9804b49w1zSpoufvo8
21bHHghJHtVfwDzzGxVltQ87CY0nPl4deBKeyUFvrNdcRuVuSDsxAQmV7O51BBVA9oqbsDcMRURZ
UTzFHEL8IkGmhrqVY1yAd9bURTPLluSxaJV02Mzvj8QdlZuIPRwB3ZZL6+OVTChSSHfSMjzI1nBv
vd2paSU4v/i+V4jpz8n06gjiYHUvqJHC7vedLAivBjODe2DF22+cHleWjGQIC6tUa2QhoIAaiO1E
GXoBpLqpcWhRLR1z1P75bEjw9pI2ObMksF2XoIpUGM0uN4lCM/0txSVxO1liEplPaXqnLIogf7tv
QaTjw6nUNUgpDPB2E0A9jycJkF1L2yt1/qwwQybI6vYya6oM2hNmDPiUIl3a32Y1ShZJr0Povnhh
9z+RpC2sd7Wi6FxPZV+yGFVduV/k4dl9sTmpSnLJrYN9rewHYpyf5mtZIrRawWuCHLq52JjppoDM
RMQXIwvBYYPs+jptIb/sVuJ9hQtyvnKp2s/QCYRKrauYTbX6q2EKBb+U99ZWsO2vl8+iq6jlyQIS
kXJbAdn4Fr/llkvNhmaxsz6etdY+asDhcTKNnVHgX0dCciETwbB3ojxkGObS7mL3hBECejWujru7
7L7yMFO4xEaVO6+ft88oFUtAmFqAYyg5Cc7aQobeEs6SaHruurVDihLxnCgnVYLSLZTosFjy1uQI
t50bDM91k2nYfeMrsrgFQMbCwGEPXcd8EL+TL8kAKO++aNf7dSKN/WaBye38uZEHfUkq0/DKK1CK
h5Zj13YIesUAEoqAGS1hPktosnyj7FbzA9Z+IoUwV0QpBBaRjI+T2PP4nrNqI3vwCSNmyWDQFpRs
lUl34BQ6F+DZhGDPMhIbfRWFUPVi7+Ij/zH61V5j8tx3/+8ael6J+o/90tddFWl5POcxqc4tGCtY
GMro4OU0hfEHcPmBXHPE0mDoydI1nIc/jbi/HG/S5XLEPhqQrl802L8KDCK6vHL7uMVz/j+CG8pA
xyefebYyn1C20amzBx1+ocb6TQyYEv8DcMIzhBZHK6qCEpFHrM0v3nZpZu2Uj9+vNMWFOzF8dMvA
LhOCRTwQJeHB8llYFPNBFmvbtWDSLaiLENVKcypM/tyoVmzdoVPj/GiEdF/F9Zel7JEL87UBG1PX
gtCliKv0GnqKoGHMiAWkDg3iWbn6gnHHu2SGKZRtL0bfzQ9auJdkLlO0dn+mq3AH9Ydp9aTNxtMk
5Z/t3Ee8IZYPeGC45m1dG41LmdtANKvNuH5W6RU97xW5+LOfhEfQJuQOy2W4sCRJLLCgTABPECKZ
6ZWiVuWqeyO2ruGZ5p5R3NhGgEO87+ISNsQ7ltNE7EnKSd6oEe7cLCW4y4nHEgG22DcanD1tHBS3
Ot3MGdx/nxCZU3Gk68I0ymVge6NGok7r+ZK3gGhUvhpUHU19K5hGjjyjRDdEVLx8SYQpgUPmJAuq
MxrOb85Fp6Woqt858K8Hb56eSR7er94Z8zcIqRUb0fkURZjj110Ttp6t9WAhlQHPKM2ag5t0B3n4
xn3wsGR7IM/UbNNe/Mvu/9PbptvXptYZYiawMpit3gvLJOxz+hAS/2ZBiBUzf4R8TPlbPwWwMG27
XX2thmEa3cHcPWMDSF7VNMdKAOBpojJdrWZj6G9UWeJ6yoA26pV0rbpEBKRH6XKh71l1CE7/bYDo
W6CcsH6+w1hfwafRU5FM4Ed1m5s1XCIrMn+ldc94XPO79BatJYCjSVl9X49J6VdppYr03vDHtgoB
9y1L01ewF3NgDozJ++0wsrVm/HILLZA7Bu4NGlGB5wxGjKOlOoS3d0WBRYhDpU7hNu2YX0aQPQHG
sIN5mNKpsbERZQiUoxyHjz/bfEaAlXy2E3Ih08nMDjl9gcuVWRkPfnFzT7nqBgyJarVkzUMpRqiE
niBzy55YAjIbEN5el9ZMmroGXrB96r9mHkCVvdGENAfOSgz7k6JiDnMNd/YoF/EhGSAaV0fuTbLa
6KBaAXohaF8UZxbXYsMJLTllw8WrhMrg4uaVNYxVH+YnC2zi3aZIjLBTryDZgQfcMmqxKXlHBEAv
78qzUoVc1xRX8xFFpxGuxOsZ0PJeiURMGbW21QBgbMqUJC20YSjOLCXEHXzcF86jPtbWWpRxxpsE
FVMLvbJeBwsCZKgijX6g0UVrmGHwKhEV/kYkbmQcvx9aYrHtBD+n2RvIj86gIBzOCR+g/jKPESzF
tAQCfOPG3SZ5PYG36Fl1OEDjVaXx+B5KWKP0IcC8lrCjj0udsjWiC0DhXErRbvt1aMRmO+TPxvMm
PAWRm9mewTKdrkrg9yYs6yAmRyly359ZyRuoMW5M49O0+pypWUWixVmnsrQuI6papiulHvhQZSZ9
guiqeqWT5vHEH5dMYb0lHTZylSzMX3gLAVIVSzO+J69+G/zDySKjlMXrFj9URH85ttoyqHmWx1CD
8YkCXPRXx648DwMS5BpbWUvndkeAh5yCEtxRq/RE+4PKHADcbbIrnL/z8BSzjoB/rwSU2nJbkXuM
HS12wmVogeb3sjjwBypM7KiIIBSOTt9y6WzETffcNZftHoFf8ihEFX6qOk2avzlck0tPfIIPpGyG
hcL3qnZwgPYeC1uRUnrlHHMdUiyxrfdhhFs2ffiW3TDSf78PlolUOYpr33YQNVqjFk/N+6AzXae/
/0w0ySsEWG7VzjoBtCFXYYIL5oYtpKEUcH8VC1fjmMG3mZ1XOTCe5zAjLRlUZ0nH1/4pS0Qh+CVu
gvkZ8mECDYcxlUPEfYhDMNag9l1AWjGbA1R2MU9ZNX2Se1YqHHHHETUEWAoKztOuHoIgzBD6CPE5
G6NJW3GGEx6cv1Hk+MqA3M7fo4XUMjIjAdmjYC8R8QZ+rR6luO0Ajtw4Gko1hZy7ySY5c5UVSKZa
8X0b0ie+DEeZWL2qux1iHxGjIBc0ucvWC3oIxNqKZn652m2gMIVVzS0hlrFH3vszenCEfO9iWOA2
lxSX3gLNVR3Cga3D5WmfNl/ggz4T4Nr3HDrgMr7ywI7S6ulF0ZgLq5bH7C1091c3DCuu6iUd75Uw
dJRLsv05bAFYav6kppH1Klp6kUsuRepnXc5+DeatQ8GvEBd/vil4lQRQ4WFG2lDFRT+qjpbd2qiN
lMjfH52qIX1ORnww+KrgpepQZanUfdeXX3ioqRV1vvgh/bQcussyGvcaILhH8mMG80QEpOyidSyH
5uGA/yAlM0D8ljrLJ7+BW3w+GvCiKptJFwoTdjvfFijVRSupMfgdJSrV5rW5FwFOQqPyZecCs4a+
IYY7PqZ0OHJ47rEpOtj8W+5NK781UOnJbURl3kVXBYmcwnvbFtdHBeOHC4Fkcj87DhjNl5bc/cIQ
B6WTetOLwNAHSyhdoIMIGdM9k9qCfW5SGHb4HjmJEwRcjiJky4sONvHfetqeXswxgOFZdvjo3wjo
/R45wafbu3IJQzXQQ6r/sWJmpTce2YUiyJoNSue0hRbUoZG/hNns+veUVpJZNfY26fkfUsJlj2om
T9Dibgj72KJd8MMwI7gQsrB4LgESojWUlN/cFYKmHaUUN9O7b7DGF9b/1zqooenjblWsxle+OpD9
hSnxVLyiLal5jH7PUl+JjmaqfYRax7Hm/jTq2jbfKJCT5H4ubQTDZwq4bfZX+MG4kFeIufzsGLGs
RKtFpNYXUU+TeI1V17G1ibIOLznfi9GMSX8C7L/gbVvayJv5oqGCM7xJ7U5mqmAhKTgsMXbWD0jY
+L30VdyByOmx0Ldi2ZIdrwyLziOrU/6rVoliGtblbAHKOoy+M9OEiRS+WHnUbUwr9ZZc7oI3Jf9l
dLos/itHdhA8OIy6Q0KdW24Iovx2Xb01BGfumnYpo7Cpr0Hll6EUnH9ZOIpcnVx1VHu6z7jmixXa
hKBzm4bFzJHakfdpGHEKAxgyodzu9qTP1N8guqlOvZrKtGExVhZtnjG6mGOfGyN1IiXJtkPvIGLR
6QVQ0fhv/TykLLocdw2Erf7lybSH1ttit7w7ISK9FibACH2whG/5Abw5Clz3cIturHP3s4us1ms0
J3emBRdS1gk67bjQMNVh0qSuo/BFD1IlJmMfuct1CQ2w+1ntQlgoIN+e+XbLb8wRn2jPBypUuXBt
E0rwwGrwTKugSlOdRwHKHwFIVphzt24jyCetuk6+ZDcd12PyZ8w/yWBURHANKzECzid9fPTEEvyz
I78SU3OIajQGkDjKIyB8gyU62/7UZoCNMEhrXgzd5fBKyt7xKxUnJCzpU8VAZ5wN1pkLaZe2lUS9
qYt0t7npj72bjQp/jfSbcMu1qrCIn2WnDAiSf8gHxFVZ3CNnxuAv9C0Noiz39X6nVWvMxvwL3Bui
ssAYNEJlaC3YFayR18ToW37J45Ovz3Hr8JvCrL7rCpYlR4rR63QJQvMksFSwvawRy5WeDx4wTBiZ
XbiKa3P8KZlhNJLJ5w375YAphi0ObBhMbeKIrhsWBcT/MeJW03UcdznaupdCFJtkITVE2y0CNcAx
IRu5kPlnWNLffOFO3ruNfkLsChYHrbMQXLZDgUrdE+8b2gHh0BcKlf3OtEOPy8C9EFhwLnZVs/jM
CXd59mmfW8jJZ8HPZcF4fbpiMhv6MABwgMWsh8B5O1JSyr9nfIVCTjLHdg7PPofZv4+oEIS2ZmTL
OZu7TSb8mcvHIy9W+vrrwzMYBMjKvQAYc+atXtnwGIiSDfO/PvWA0cW/4Bbyh6bKamsCtFWE0Gar
NUji9kL3eryA561tfvXI9mE/3/38ZIWHWgaiIGAweoxMcEJ57AS4dwzsPULHIwKfDk8S6TlA8hw5
uuqXhl476rP54LSvs1cIunBqdzE7+QvZNejB2WyH1IFvk+T05e98s2G4dapPiCLiDK0klB+uk2KV
sRL2RpWPKsovpHEozCXZ3yRC6vx11ECKvceqtB/+vHEFGCXex6SAvmx1gu+xzFGhsfqP9DU7YYzz
1XiBgQxdSh+Bduc/xUrvwFxgq+qbMFXm8QhEsY2lSCTADuxdQjxVAaji0QZ5Qz3Esq0na0LkkG80
6pywxQk6q6l/A5iQxqV1JG3VAQ2k/GPya4Tc+CkAFRSrAyj6eY8Kf2ZT4jbtOWJAoW2oNCt5doXw
QYrCKhIZlz3TwxUXtjwu6qgXSybF/QbP2OcMBl1LPeezGqlOAarXfiazENyp9Pw/kWybQErUDm5I
7vAmK2TeUC3/HAIHf/cq1ssrSAzCVtwgb4O3dgWadlp1Hjiwxh86jHvGyBjSYu3ay5swsnwOdL0N
q5ME2/BE4CMelV9hWxH35wPQ7N5F5crVx4uRr4mqPazPSF55YVXclrTcx71tKIJxyZK+WVrWucRp
quwNywjqtD1hwuwSNJ59+BnRePNIH5Vs9vFCzhSAEr7F1GIGKo+wY+jJdaMhb82EncK5q3kBHBDR
TWG5JxGm6OFvvkTg6N+pIt4nF6OgCInAs2fXzStMOyvZU2fgneKkfvdHcWU+CaY9M6TJFkSGTIJE
a4kj7XdxH8kg3cqcRevepp4F02clF+pl6/WHITlC/5YHU8H38xTnX+FYsZP06HlsQiOkV9aMVBO1
rKuKgKAAl5JWQijqff1lfO8GLJQeC1gSwD0E5TzYHBs94TzGZtUQ598sbc0jK5Ta8OL9nmUEti9e
ho55g4zYuIzF82hKDQtYB5wRgwfGawBi2ip2D0HU2Ra6GaKKV0gcCyI64rMRbIrdsS9662GVeaSP
ugZk+OO3gBq0XYUnZanIEnLmQspDmBPc0ofvgLATJRxtKD9Yz2qn7W8w8v2LDnIIjhI2oPuMXl6I
lzRKgmb7PBT00Ol97qsm2LNANQcjh8RZ1ZRfBBaKcbtf3YvYHPgi68oNUMNMJWNupPINMRY7IS5f
fc40yZyr11KOzkfix9LHIfjvX57gggt4KU2HkKGeU9xHrLrBV20xEwIcbzd8895qd3HT1HgMeDVQ
74EYiJhHLG1sPLnzzzxwq9b2esEkMU5B/1DOMdo/WH19en1zKzUwKCESN8PQq/S3Qjody9e+ORJK
07KydGsRbibvHj+eJVj5j7g39tRivlNQbsUdAmeOOArUvZlyWk2ogh3NCPO6tbQhxBogGnMuH6Ik
e8XnWzXhRJwQh7I1DoQVeYa6Di0lfJAWVICIjGeEU1s/z3AUbZuyKZLmyON2TK4sJ51+hnG96O1P
gjL1diY1BuAc//cfAnMXMb5by41sFKA7hZ/LTk9SpvVUzEHSVw3jZ9JN/gg3Iv3QAZSN3KDgy+vm
T7Bk+GEl66oSxewe412ojVt1nmaAcaI9nHE4FJseS/cS/PP2vW4qPQnLbJZpLGkVU3pIQB7ZDIHM
qUjAOBSL/7a73o3JWEpm+yeYAqkr04VHA/nOHGe9K1kzgI9Ynm6GyJzRwMRqEeuf/8yJCVrZn4pU
L5q5futMq/2yBwEvsBfPYS2eQymXQBHEH8WUotlEF91xLPh3th9DOrO9iY6O2/R6PDRT597UhSbs
S0s+z2yTLhO34X4iVr1A3X4mjVYzm/wG3Yh/SiVoeCPRW+6k5Dem9zWj4DJMdTdKsk5fHlYh1ud6
rsxy1ZXdrNculze+CZ+2aSZlZjfsb8hPCDCmDJCA95SqU4hLvkIWGmSnjyao3P4Ye0jMlvusqj+r
ncdJIPpcloics3fekamEu0lL4SmeEsp4qV+NYDPjo+wlSXBhJAenX7pk+z8bXZchjLXwKO+LEx4e
isRa8rkCp30+AHRc7XS6ISp37R0qXJXJKQ39PrbjB/FfWVShFGw+SoyEFkcXVUqpMSESH6F38Zv4
9S1nLxAQZ+v3htoLhwvrCWTaz6EWs/DCHlF3RY86gzOkLGWCTOgOr59xxvkANEbkSHWKkgXuwnVT
y35h9s58IzUC67Z4dimmHWN+BhGRwxFfSePD3n8L7CgkwH6Z3G3IuftLU6agjrLRqrb0Oz6h8eBn
cFP61+GGbaXcLHpqcoczJYx8maNRCrfOe8qIZHaO+HkynvedZ957oDGRuqDKiwySfns5bfNn3Hc3
h4wUjWXTOKzK4kv/5cuPjBnxIv3RO1QUHRz4oXk/zUINNtXLMNxzLTNOU9zyTJmMKejvwC6SqZq3
KWQLSh8ZWhjRzNtg6//hkx9sMW8v/QYmY9HVUNpiLuc7MUW6y6/8fTczq+H7Nmj2G5Pt4FvYJ7UB
ryRbml6VaDU8RRwlM/1+Q4GdAYaa1etQeIBErd8fYKtqByH6ClT4fpxafgJ+IFlxyn1Xul/hWa9h
12BgefX8sm6PXFThcVcuns/8wPTfEV4LrCdA7Rs73KdKeTGWdslrZ10JFi3cGUjwpyuo6zXXTSxQ
p0iBVjnK9bOQl69IDOic/TNjIGIHYlwJAr73OGHqkLh2owY2dWz5EuAGAXBQgpbZ4G82bXzZr9Yo
ZG197ULdmubGzrCld3kcU7yd2SbgE103vcOWD/2Qzj11DHnlp7QNddhGXcVK2KhSuIstE3ggfVzG
FCgrI0HNrIMiyfqkliqrn4RT2j/CNw7OooTF3hObX63f0ciFUPUwi5+0hwQvgsMvLQSJ9zgSLH9i
3BXFitRvBui+5/5LhqGnJ1KQ6DNm/WdQkd4SApx1FHVP7dokM7wlWHGLiLBRY0Z6p76sPA3zLOiW
G1T3a2HywDdyNzmMIqLAfEHfAdjgc/YcrP2ifA2lVVadDpZcFcW4l3TDMxruL2Vgp2G2RNco1HQb
XMwM9qfjXRGfmkEQXUVShCeFyNhaobcgIPMrCEhPJFOSeNucg2RO9UAgS2RxcDUDdjk2QyOlDUiT
G+gMnytaGynblXmNbwN0GMd0c3apGu/NuKyQof64TwDvQeNbuI7AMMR4cpcz6NlGJPlZcW0HqTY0
+XFFdnC7OjfpC97yRe2Ycj6FVIwEPnGmJ9OYNGeI/x2mlHshsiBDrvdyNGZAUU6Yi7z5GRgZayLn
ybR5B/YLU7fUDMaqnE5OFCb0gJXyHRwYVPtxBX/yQjFC28c8e5UtsT+xcEewxPzYBERFYwzXrmq5
hzdvW9w5nBvTMJnBnYn+0qwAKfET6w9j3PLJ1Z/vVM8Ha8lP16KOeC2GzdkQbadxwRWevQRK1MIn
TbYA4drucfNabH8DNQl1vCb+zFwOXxpnWqJ66i5bVgZEGy2Etqd8grjfTM8JL4oiI0dVlSYWinf7
xASj9JhJOkS8/HtFEE4pX5PzqUHG/+sCb9Y2Gks0/6dUJGevTXbPvenxwEdXYa161MMVT9ViNE9T
iwKWKtFAJGGoS8/4QBBVPyx/PArwsKzwdE2zZRxrVnPwwYx/DWmN32AgGbYPai62gLVDpswO6+cm
dPykSjsf07giVI8eJWNoyKq3krUWs8tr70TiaPtSm7cFEoKzc1o2mTUa5lT0xnyr8ZBV+SVCj4tp
CGxlBHiMV+CvX7RATHaQqE3CJWEC5GtVVxe6oQNUHqZbEMsLP0oIGuPaa5D5ROx8HtF34XsuIFmQ
Zo3jhZOH3507+dL/PiT5CspHUXe2op0gEVjh+T0L4OUlx2E4SB/kQ9mjsydcFAihVSk7gxu30wml
JazyDBV7QHDePPwSU9qb0q/wqzQzbTscXfPz2nC6PpPqWic0NAhUu8fSChs7vNP3DwGAYje9UB/R
SdinkmWqQRyobF4qYgj7qxtuwBkUFVChm++MaZjJwGvWlYldnr0mOtbK4yb+onqu597/xYDjV5BM
jEyV4BHgaINKkJClR+fxe5hMMaMd/nQGCyTjvrAXFg92XfIQIo9NNKiJSIGcnefrAvDuZp1bVvE4
+kWl9moKXkv+kV+yW6bZWBiL5vw7ymbN5vHUNtw36AklZomNondWIhPQR8D1gkb+sXBuMSSD6fkQ
ciUWwKojOpw51mgngGTRIXOd1rVt7tLu0zIbIG304Zz+03v9h8/Zlyi8j0o/sWtUQwkZvaMh4Qa4
1NtJyl6prRpKt1z2BdrS9K+825ZpqGbSD5WWeMyzy3EjOZ9EuuXblbEeafz1ojVEdEJBKDJZ0AQl
6tqCESzq700xD69M+lkvxswOixcgeqjBUbmPpADWYEM2u4u7WBchIRU3OdH90iHnYWrPiNDysEtT
v+llPQ/EgU3Ak7olhd1S9B0lbzP+GIBL6l0IlCRGuushiyGIW8fkDNIsaEkY7dc5KGAl1meqNOBU
nVvyYKAK98fDAsGkwYHsz3pqDz/1u4sduV2qLzr42jUWV5RsW63GRgyucg/n6BH06/D9V/8droTO
PPNtyI/GBBy7by7l3Zq/wLda0ro6XyJnjXp5OwnqwkdXZsqK8LlqGp1N4yCRYoyzDe47LAF9fpv6
IHP4LITEVB1yLKMPu/Ur5yK2nPgNTKr4QUqx5/BQIsbE+MaRRCZuTxQxhBlA8bQGmYEp6VDzVftI
duhTPNYqXWozGV6u0IWAStGfIDdYk2BNdzkMb2wQP19q/NcCRWYdiooa1hGt2wwTZAQJAO2v4F00
QAM351IXd5c1JJ1q2XhEWKB5y/DeaL3mv0IL5hGdK/heA5gkL9zDkWNcZiqEKR2itviQneXtFi00
MEE7iK98TO/GMca3kREQplXhU3GYCEvDXEJ4mGA9wI2lMZz+XeWRNWOMKiQp8nXoQmBCMN6qqKse
+s45VeyykzAn+q5cKcN3tKPGgapNQcr/Wgq85pMdbf/fgqDTKGwHllkzMlWZB0WDYhWVj8Og7wht
/PhpG9owZypVlMVfwU8inBAt/pgNeFx6ZTlKqB4690lSNr8IlTUjnGZIBphEMXrswBQxog4fijys
ReLa0wJ7Vl9aR4Dbf6O1rRebR9qoC7dGTCiQmplhYCN+L2EhKqDv30cUuNyhAr3W3lI0Q00b4tBk
fjjVEfASQWj3Hh4xo1zKl6MNoDo+Dlh4topbL0bn32EySzMWTx2N4RWdIMAWYSgx7fE0/BemsAU+
EILO5wJMktrjRYxHpH+VIag+8Wy4gjUIrlfdNT1QpR7cgghtN7CxkDfa9N92tlzTkxpkme8QqTCN
0QzpA1H/FpGpKvkQlOzMhbFXW6x49U7ImkHmk7rP5cpw+sFyw0cjY3Pm9usqBbjyfYXSkSvVw/G8
ohpa9GkVEgXYvtbTq+Oe3B5IQVG7WA+GE+Lqqg97HkOF5g/zDGckbPZMjV3Wa+eGCSizq6y7JDE9
vmUo70AA1ytQOacQ13b1lPstIAI4QZwlWEcjyJsB7ToKkBW7HgbC0LuzetZaSNTtikO2q/KGjeWg
aKnXVXOz9PudMeo4vHsrYEm8HwriPzxvIrM46o7ONngS83uY9FjYbPjIjZHQ+j+YlNb7W4w4rsDv
L6Q5vI0rQbTYVpW5vC27oggEydDuBnvIcaf7R5uJHEzBldDrgDCSBUZaQfEUBkYmiQNBj6zogisU
vH//Pu+VhLqUpGjf52lUyyVSKY0aNq87wvR6kfmt4gY6JOuMfef90aXHMGdldxbQTK8wQU7cUwns
WZn5n9mlvZFGJ93YVNjwpZCgFQEg9jLAU0itqvcOr17rStA3OvqJx2wBwHyl2lGdr+P0474dVdzc
igUvzgH7rjkVqf2QyD0ldtEXyDT8uPeKKy7TXExco376yheh4Ip9uwCsSdPp3O2yUdy6LHga9vAj
xIYg77fF4/h/BT7l0pCSH/8A452/OxwfJCsYLfB9Ug45aDmXE6dvVGC6FkK15nKYTjQ2/haGdP1u
VNBkF+cVYlVIKTEzGtvH2dr8Kro+2qwJZYXqbbSgz08vLVqN8DP63Q8vVsPp2XSKJWi+Mdevz7eb
e4I9OTIlfDqCZEdiTSr/IJZF7aqxHTprQ5DAfDdyBY+KlY8OW7GDD7wiksTEmkTvmChtCpZJ38Mi
/+wboP5fO4E6Hw888JkdrSyc3IRfMiTHoyyHFINo7E3m1duCH7FO7Jh7G4vUnqQWI9/CQMTuYnrM
bwMtFLs5pKALIkT0LC/pKsUZo4VftW6GMhnWY6lrlnHENtxSLGaT8Fd65wCZBBlstzpqlDgoF7D1
k7ZXr2s4n3/Tlzuj/8t3tvdRyntOLJdZ7NKvgGrk88bjVTt1q8B5oL/Mgh+6TDvAg6mJs8s1jnOY
B5sfSbA9MLQcnKOWK5m3h4Ksyq0/U9mX6HF4Nz10PE3ssgdeP1xwqveu6F66zsvgyTknHOprDklP
dqT+YimIJlTSmY7e9zA4HUUlixiFsNdMDBy+UMxWb+vsd1r+z1UG/k60elzzXT06D3tD4T3vpPnh
sK7q6HKUi7xT4nw8X9JB3oEtVaNSjmbz61JtZsQOzJ7O2tWyRMZ88pRFgs5o36hBWm8StP50NKux
KP9psPR8O48KWYqzlVieewCf1cuK05XrakTEi41npnrzp4P3JKrK+KvkKa3pa2+dV+Zah9iHXem0
d7H0Gb7bRTJHOu6KA+5OO502f+jf/gfWa2a2XnKWOGCBFITgjV5xJ5pSQBq+4kd6QZBKIHs04wpO
PSb4Qr0mvcVluzxaJgVYRtoe8fUFZUP0mTCoQJeRgi0VGLWPKyR6R/CCs6TZreUu1UGqZf8IKzuQ
IBw0dtpyBNZjhYvcaVdSGs11j4ZynVgezcdw4EYvmRvRxppU4/o2+XY/LwqTIQzKxHtZ+tLVJUW6
mtSY7sZFQm36u9af02Y1YcQVx2SPacDcbwT1KXP6t+AuGhOLYq+hXpErLu7vYdAzVwxU9lHIMFJe
5Fj36kjIUlMY9+2YNClW5UvCtyRPkEGwqtEfaRP52NNmy2M0/8Tb87AEO63gamAUMNS+uFNkYVxt
HO22uaz1B+Moa12gIRahIw3Ce6a09v3+9qwpqmbFQrDwDzYvQzogF9jdyWoFinPR393yN58mW+Ie
WF8rMl8qwFxlGKmFdOyMPSfGUvG8KXgVS9DwK/HQ+Lre/ZqFiG1SWMb1BD2Dd8x+DMTNPCuFsVTp
NsRuBnWwl0jTy0uvReoDptLLVtMxt6KklFo4MWsd1Ut5IaHn2mgorn+GInVO1SsM4H6pgaZNAjQd
ojgi2sbFs5jz6HxO00vnUVvcaiEl8vjv8LNCJBsoMXMMNHdTK9NRCxYtLZKYD0nJb5hHRjTzDK10
q/xKeUFhtOkSplEWWR1cAXIJS8HyZLTJg5MytvlwL8eeKr5ytSJlYI69Qjkdw1AgCl4On7wDkeTu
T5whGn8ncv6GAYeVBJJPR8EaWA5nttb70H6CdyhCVSfpwmHjEP8HJFzPnoSME+BqSWq3Ci/sch8z
pLAcu7zSJe0rRoEhT+SA6GMYe960SjZxF8zn+QF44TG7AL917BPsY7W6+doABDvjTLA1wjqNU5rf
hBXkb6sTHbcrjMlQmKVMMmNC6AR+OVPmq5Rgkpv5ccZOJJHXe43mu4WVSXy+30xdmS0L3zEOXRTO
zMVGFtwJXjlsw9FKrjLYcb0VwIRTiRG5Ld/Jg0PGnafi8kyTWOKyGTZWObBrqXkg8xv02eH+ss+j
yEvD1iMU42U/UFdefTcZIgJiYPSajtQcvuF21pUm37jPZmdVdA3DqkuTwWioRFvstLVstqasBH0o
KmDHV/b4yQ3NAkYqrjzRqd4/v9o+AlNTpHcLxT8qZrh8wvC5ougSyzVN3Ae7IiDNbH2BLPSK9gEg
kvRFtU6b0WCrYepD1QUipstE1qjAZSZc2CbRQtkQ+cm7XthbErM+MCvpnY6gT12c6w5ACxoFwwBI
luGx9/fGHuAXv/wX+Hy6oaQ/SCs2xWfJUe808MKxlzW2wMPfOx5+I1UqZ2Xs+akYiDhux7LyRN/+
XSj3836ndznsfYietCk6Mgagd8WYeUO2DTexbt0sABrthGMyrpev3vT8h1YQQzpMpWzEBSDX4/Kd
vDSJSJ5KGRfhGUdS9sRNiHKRSfKNEMlgO3HG4r82zzTKHI4i0UGjXLg0ehysaOjbg7jf4moU1AeW
T/vtE91rg13rGZybtgI0CzZgIKLwlS0qojvj8nRcY3dSbeKhA0PK/19i/22E2B3dUAq/dAEfc6RD
mRV4hc8HRop3KvJkX4Gn+dIlzYtHVT5VQYjwuuaRTuIDj5p9ZwNLKXIc1IolVnzz3hlS+8Yrya5t
ljJK6VJAz45OfjCl3gVIOk6wHLQ+yGOgNoJDxEWcAWW3Bv4srdMFUfKOCmxyL/3rjdqz8vGlF6X8
T2OzGttAko3bMQXn/w/gyxtmKxme3DLG/ezlT1g3KMDwn+kVGaFtjHE/NGH1YJEPwRQptwm3C6/0
xr7j7wQhZhsJajgDg6+Mn3NLMRq7qgcXUH/wR6VEg/cWaHbGKqfqlzd7GThf4/OO7W9iepMbNCc6
R0ptG6dTDuUtgSRzKEIhYZ6OpxBWnGM5egbGvYEHbJfYIuhoO2x6Om3GvBFizsnpgO9BbdoMLuUA
UYSgaptct0bmmjCWe/W4Bx5QyZN0pbYHcxiXzZE1LnpvQgKHUT3bo40TaDwE0QOStZdCuERP3EAF
44DDRMAeltJvI8+RgPWGAQI69svvWSm68hH1oLtw7T7QOmLTLkvTDiGo5P7cyYXZmeyV0uteVmiT
ToqERwnW8Sux+80IrGOgcV07X3+fjhdYQr8PJZts1OmfLcMuJf/JvANfAVEAyNQJvnHFn5nPcF0d
oog5ZjerOrV2eZY1NFiEC3CJPR8QEfOZfiWCx5SLBhn7n4Mh1zjvkjwPCQ6w6DuxLIMDQFFM1/zX
TkloqZQXFTaMztGjTNlKmhA8ugeNvufqZqW+7bWXk3syEPnjLVYDwjfMXaDyYlf363sIcHnx4qgf
LcvXNIE5knTGiWPnFqyNTcY53bt6XDkW6gt7piXHPSHkjPP+EDLoov64qqvenvC63ujqIbalwjDR
VpxbSO41/zooyJY6uS9vBOvyiALQpBzQfuq3udBu9JYBpA8Q/dsOCgMmBaS622lKqCz1N6+OZFsq
KNPKFBfnEnkh1awaCrCNlMkZjp7P2yMgpNbAwOPCMcI1gY4w2FPnyQJSdA2bFGEmQSUBDXdXiU2Z
+A93SuDIhi45Kv5HhyQ1DRoUrEMhwazCKclzMuELpovvH6bI1Ib1ZwNPZKfh2NigxZh0//pqNpXV
AGb+lkrUQVLxSI4jPCUhHwpts5xD2VWfZaC5XHmjjZbfx5bU2zFr1vtu8ynsjeGtzm9SmLJrkQ1U
fcPLdJrJiCnMHv4VLU0NNVAbkiYQTeiXM3HYKZINL1r3YkO0Cu9DhzPU9qMtR1McgJVefPmQjxXI
D57BA3dwBQD1qlIifOhrbUYucfQSfuI2CaGLzqtJPB1sFrPSZf+bdFOZSVLfPibiLJJW1V0DOZYs
JuZxnGgm51XoTVxdTbwqzy26WPH5gNUayNH89aOY8LcRrSi8kRkls72nlFsGawvDTx4enj8LLCqE
fgBmaV/9EstHOLqqv7dkDny7XtyvAwZZpkd0IIxHPZOjL8mqmYW2BDYLClWKSdq5A8+Ym/bgwyX9
WajcDAbx5FEeOlHs6odKQor3PhEtIVfuhoTU0GJnKKEb4XX0T9FJDH0y3mSlH9llx95eBCnNTTmm
3sZeVg4kDdm2S1qFfNjgMDH1nX1vZw6WsirZhtKnqWAbA5kaAN81Q0JD56cP500DXrIhap60b0V2
PPdmvKJlDHaSPTPe9DzSxIVU5qJRLseWElt9RikLm50bq4kMZK/DMAMGPKT7RRwG2Q/vsyyNhIYo
Th5c39eVO/P3DYX9WYrv8nz2fYjs0ttKxzgVyLgcb1Na+7Msu5BDNIiTzFA/POnc1R+eDv8o16XM
YT8QU7AOVzdFPDS6RevE+nwTlqQS4Ffgg4gGJChUg5fLXzGNtiGcbEZNnDF0TkLnSPfJveLHqeZf
5tAlxh8tLeKRWr9UmbUG4w9uGtDUOy8nFUp4xnkAwln5wyl0LdBoWUgriwvz0AB4r9FOJCl/hEQU
WraChXFBLhQX4/WYI5azH4zofmUUJMueZ/bZiRJ6fJ3MqMc2+4yl/Fi1sgPNBr4RcvBAJciiCuJB
5bHRP5bREftemVG7uV4/1UIbievG0teLHAQuXddX0sHXgIvWXFn79pyI126niVD/pHt3tdndX79T
AyC7iThWEMmV++MDMJx5Prj3CBgGBMAIKScpMk5d6wK+zBlLjtK5IrqWv98MxDtZqfYm7u4gQMd4
+H16MzP0ISIuMKTxpHfI4RcLHo8Vg26pwqT9SDJDK5kPIVtIMJogE+tlCvhtM0DgJ56146oHsvkG
z+nvzFdOxrlnCqYNi4GkmnrTn2ueJTf8/sK/m7jn2JRhuVRQoMxh6XctE1tjqjyXoAHuuSq17byN
Uj3pA2gVqDyYyhXKIYdTqJd4nvC0fupv+cUpxYuo6UZxPp2HA1gxCPwI28l/lzFugQk/CjAEr27k
S5fb8ORG9ijF96LZVphvAQiI2WIIrit2dCdBdnrfH9NSG2rUnB3tiigawaCnteJpX5Ug7EMnuts6
miULAW6vTKl/11+aJ71wsyeH1ro9UiuxOHBSfTGf2mrRVfdsdCHEm2eBqtRnZq4rGusA0vz+hDec
KJs+yIuVsXs1Dittiqoi42MvPvsH/0gXshQRxMmgXsRh5/2c0EOkIS9F2ug4fCokEwpsr/6ys5x5
JStUYZQkKFzpZ7KFYjFgmJQ277qS2jKw92n2YioTdqTRuW7byt2bTXd3yNnBcqTg8JjoVDaWxuV5
cJssngcuYfpG4W6LXBSiaqNhiFbpLU9CdSlCbLZuvJ06qteuLhTQweq1r7R5H/3kRb/MExiNrVFn
GjmaIny2rgX5R1Vz5/7yHf3ff/rOyST0WMhE1+YeCxLVQ+LIu3sgrps/00n5Ao3tuadRRIMLi+hM
fNPsPAJzniEu+OB4ltcDa+lyci88bRAJzq2swdDGb8gEcQazE2Y3Ut0rNOrEDgQyMphd7NbQO8im
8x+puTq2Ju/Q9p7R1gkpIuVTlOES9Sa6tbKOYqFmFRikBcpXjM7mC4VemZVHGlKxtdqLmlUW5qyn
OtLMyTI14bVyDhwWC2MJk8msmYhZfkqDZj7lAVOT22wRYNLIFRbJRhj/XvwMkVaT/xq8pY/IX7uK
zzBeruA4MFpjOVetVJdLQ19tG94nuaRCyNXGG/7s08MbRpv48FW+9eS6pRGc5mgFbUWMphhmuP5j
l/L7/eOFPuwie+b1NIZCFgEl2/lx65eBStmrD4/vv8y27xqz+j6yVBPMtHi+1VEoKXt3GxUqgliN
5Yl7uscMaEXKq4yyNL4XDNIJ47+uMw/XiErveYv0NbST2hViVrwAyQxSdft9PEijltwjNEiOCDRC
76vpjPubL3HVl/DGp/J+5CPB9H0W7s+lrcNm0voIm2wYp0paOcRankdmCYoiW35TsLh+UitLDoji
IP255DEZhlXaaich/4xf4IRQZXt0ZJYfTdSHNHfBUSEeT1Oz4LlwTx4BKCy8uFJkbVdKhd320nDx
5M9oHSQkAdKYckIF3fLgiR96LqkFyYNMKzKN7yicWO05rnuzXliklOpNslt0hFpUsSmkVd8WMsla
TtZE1w5BAv30C7Fn32cPMp+gfQmrtA6WuaPISjNctwwTUpwH+FfEu6mMORdgduRkgCKqBH+jw5lo
CHOGwgdDPpy4AOBtOyqgZh4OlLixTajoHDP5BDVrSc19WWuIj6FJg0aEEYwKImiDiJE9vE3MJITy
JObg9xrVt37XGBUfDYGUWZQ9A7LGHI+rHMPBuOyxkNQ08bJSqOYVanhK552cWlkZ14/Ve2lH3bM5
TzUPseyoN0WgUGEUxnj71hfaOpJsOtRi7wzRU8b2D6ZMCXBIsKnCyEDo1dkaMLyWKQcfDjVkU4Xh
H4cMxxEBzS5VHQd0zHAVUWRRXKR/Vj6Qp8NKtrUliW6eeU+QxGBFhwZAFuU7QT+ZvEZODYzS19AU
fyEy/O/CJrmqZ/7UpX2ykR4dLC8V2AlB5CPG7aArSt22reXXqgpxB6iSq4HDMu0upnntQ9w2yT3u
7NzT1pwMYlJiW0v3FhPvii1AoLaGfs/WpE7BW6ym6OC90sy5ugQ6mVfKZw3olvhpYq7wTIPCSjHk
u4RjwV9Uz7oxVsuzIIr/z8Dm9Juf+MYzDr4IVdPuiBHSwj0RLUHg9RUIZs9mvxT3v2oUjZKbotkq
cByweT6ldK6gko/ZYJ/zNwRUXxVrkqe9lFxP+wkALV0RsE0Ms1MTz/stG3T3CX9Wthm1Ep/IvJls
68RZHZsKWVs+kwOaXXVFO+qsAYOT2FGGrsguHyRMUkNWRhoS9kuUKLOYQYXzT5qnHD7qk/rA8x9O
iCEAD/WNWECJmnqDxeog6SCv7jVRjnC1vDDlc69CDEBbVG0wFVEdY+k9Xbh5pcLL7DTLXfSUU8if
2iab/xWncC/luUlZt/qDQT4PgTztYQ7DS8+0DFaHj58TxNfxmltMFz9npJ2KGDmWh/WHOYK07TaO
C5IZEufB17ErDtowMekN+ZiwdqamoEoDtQrwnABtbLOudgGiJwuKsLwqimFba/ujYJg+89DIK9+I
cTA5z3/dS1L43KkDAwua+GqKrk4yQMPkMjTbE0+CL4+lG6DJiTI+mho3j7cxCfpsdaJUSnVS5BIR
LlWmwgIBNKFMJOS/2T8pdwwqxWfG11iHihd4WGewbKrZY5BAw+lwBXF3gv4bc571FQc0mjg5O0DG
+NCHh/EdKi/fk2lOHR2X3zukt2Imf8ygEwazqsPOzC5CZ2u8wbSS+Fzff43Su9+ycn5ciybAYjL/
TSlWzhwfyFxWruHSLrLWGP9SBFGjDaS2WbnM7Sk49CT5eHNyQyEcREOLpe0Ec61IOXA3R6AeoXC6
TbKfsWeKHncvRFb9CmRqQpmhuNfKUpb/EE6bjGkjYWwfr0ltBkDKHXn1J6GOLUPsz3TM/rjnOOOr
Rr/iVVmM74FvW+mGIG0VVQd9vhU8OyWQMBESe5zI4fmH4yjPQDXKaytSfRSDf6Fw+2LRXKy5YOpg
/VyWejKdtYIN3kpoxJ0Fd3J1hKlTKGMLtgnYmjxDhdpNhXYcF009Tyd9635GrN0+d10cHTnqcNUA
bMs6uMcQyXZg5MDvYG9PuGhSSAexx1QAa/fFQPUHsLeERsSsW2mfQdqJY1QboAp3rAOzeY9x7A/O
TxfmZ3wq1xSLeTjeOOyYPOzLNor5KyLgpX5yYlX6mYRksv4RA+wigBtBZaChfRc14z6k5L/g/HoH
cfxe77KitX9fNZFeUnbCWycMP8O9QkKSbhgxAs6GnipJIC9xSrRV1Sbr/pSIEE5eQ92azPgBPITv
gnCC/r6MjXoLMjPS3yI+28ML2f+JNIgzgwFLx0I9OqEnL41adSMWZeHNjJyd907nO1icARoatqY6
2Tzxrn7NDAfj5o2e5UViWRricfs3VObElQcF3VSNvQ02sZKhp7q6Y3KPOcxT7gosVvUo/VqeluYT
3XLB1RhFGpBQjSF/b+3Esju8YzFbyNvW5I4Ct4y0YqYU5RQTnQhtaXjjlaDT6J5UB7osz8zFEUQw
SaSZ1pYUOa3OMRADbiMv0VFLWCzS/0/dhHTeZwPD+lIP5ZRNzjcN/hGnPV2mXSrf4D3TJjCShU44
Ch83dfsc0i7+ti9EX0a6jLbN1FSBMGX5s90flM37+hP+cMVImzSXF7DD1V//+Fpbby36zGFOs3mS
UDGKnb+uaTLWodOwZoQWEWwGB9XT+aVxPh3lBdU+8FPAp9Rh7MnqvbH+/E1lBr/idDqRGdTTgMk7
Frp3NItkGTsJLfW+4ugjmCG2DQx1JsY+RNYGbHl3Qv9je6FjKewvcKnm6YyY1H4W1WCK03NIiTao
pnM4L5GcIx5ENH7HhCilWpMZXax+Dk3Lwhkq0yCA6a+L4hz4ZyJ2TKVzKrWI1SmvhjJgkA0DGpEY
VoSOBRtT9DHWzuASBCQjxvQDrng0kfDkdhTiSKXxW7h9Dd3qLLHbxVoWNQTwm3skSimTBE3Tb9zQ
5VKZPfoyuXezRNu8QTrSYgMiLGXXS97dRdJR8AP7XTxlKBs2SfscBv/lq4pgH0J5yjnGxQSbTNpu
eWl7p3dEFict36I9Gj5OoJn9Jl0zcQ16yu6vK22HQs8FZvFYGjgt+qHA1z2IilRbvTt1R+7v4qiw
ylAbFiUU/A8+0iCOjN90BNVYhxXTdoBUC5u53FDimm9dhtKTrJT8DsRNYwXmsTIUE6pSRqZbi2PX
JuJexMhmCczHQzLPwjxL3nHTDi9TXhAulbiHRgIuI+iY+BTuMP0z1lDFbdyT0sZWfLULr7kRuzsn
YWoNJXwYHp8gV1oc+HKVZkHLlmwL/ADiiiL+AXYP/1FCE2YyzmQmKO+n0MJPx8bOnSknb39wNs2P
UkvuJbMqVVhuiNdeZ6aunV9DH0sAEuTRFQ3fzNEf6S2RWFZj5gmwbny2+YMJrIlGjO57svO7ZANc
em7G+6EhOzU2ww4wVc66GskiV4OvdRylnC4+kQgpRSJnTgFtQk4RcwdaoeG4UG9SAyqU4bFIPRGV
LuNRfwcfAd5ZKPYrCvvCpRJI629z4vD1AJfMxkaqkMLuxyFyy+Wc84NAe1eM0mLsQ7loBm4BQ3ms
2t8uKNydiOXjlpyH/ehJ9zMtQKhEyj1x8PG0srYz8Ot90uUwZfsLkA40lXBFPhS/6q14oYIPU6Iy
4BwX/Q6lb6tHxfS/4hw+7UNghjK8+X2pDCFwj12B8AbOlOlLlabr5/2DlHpVdYeAgk+ayodi9DZx
quOWcA/LTt2RjWhGhuTMdrhNM+aHdXZlRhiQlVo7l55w9TC5owJNav31USAo5ccDnntGZADMlJeb
hbSaAynLKda46gcJjUNhnT1L0R0KASpvu+r4exLESxV6ApW5M8lPj4ksy4trUZurFPrDi7uH5nGF
Soiky5Cf4yurpqG0juqNWiOP8dKPawOC5+hqt4wVsuD24ryFF4QNhvqiC6k71YHhlx75lXxHZAgI
oIhPWliLniLbHkXXH0K5Hbj5XSI6qbnPSaL1QmDEq8u6tUVf+sO9BVBz0X5DERL0Tf5DXQqN84gz
kX4S6HRjxDAkSVKPWXO3hSxYhnAsRjnEqI57PrSbMXpVR6X2JLu7l2iYvtf+VdS9ED0xDs0x8kCy
5wJvlPLGa5kN/aOoakzDporFSkHsgYbGUjRlc3ElnuMxFVDcUYhfCChnorCXydJK7N46b/WIOFOr
+DF3RHZqxu9Lj64aLghzDvDK6K5y+OMouKl2QUK91lZaQpM3HYdXKK7ApIosRw0kKIHvIcD/O4mI
CZrd/Lla2klbsndfKf7oPI8l2/9n8MsXt/Lj1eo7JQgHdTnUYa80vqSeKg0R+9l0IrZbhvIlOyTv
xlOzVsC8bzFTaOIQoUlRkCqmnKs/xAv0cFRfvs1KsA2oZPmullLC2T1/jcRcIlEUB/JCSU+qySTj
QqWarMg5dY3PmbEa5XlBlbQDn/4c39p2e/nFo2isGWZm8typiieangYjxzZFbqQANNHj4eRGWjyT
0lIYMLmIf0rl5YPJkF5nFxmWWz9oLWBZElP0F2JkOj4tHRng9r1gLK5fv+sWEYP1wA9OR/hIpFQw
R/9P5f6yCpfcZjzoygoID/ndPRYb4CTl587tk46yJF8nE94J/lmhAq6PsyivO3WqTQxrPlNL1v5e
xBSAU53e4GE6JDoTQjQg5d5s7DS4Vms19CzfGUbPUqtBZdyolSBuP42SSx/eNxFepn7waQcyxhQx
ZqL4tq+I8a4MpuW9yz4hMDlI2FwwGR+qsQTlFHGaFhzGJcXsWIPkQ3Bap3uW4UtM5pz8Qf5DVxJP
EPX0yRj6OZxHtmqTASbzQ8DznkFSDSsFm82A6j54THeSpZuyRnEYcQkAeQkL40T8Zu3a0sYd/qqz
q3f5BqBjfUnhzkOqNYWmW4/EuE0WqFa41kQ+XzZG5ifzUghE+2J5O/yEG8BOzs+jtXwhwphH2fjJ
DJHkw4uS4DYUUo4d/QdZnpbPUV2Ehq86Lt/MQtuTQNXypeJhzcxm3YDYwJmcf9h0kW3Uh/fyZHi6
+jz6ZMrnU/2Mnnvm6ze806nDQCtNHbjIP/CBB2/1lgRsZqs4g0VBGdHKjeg3GHfCnGhn5A9l5NkI
QAYkfZsq6ngXmO1i+ul91ayHiED0OTmavMr5nldrodCWyWnOxvAwv4tCH2MeB2WI6V7Mnelr8lr8
nl27lSizgGt0mHB6VoB7Q9h5Ryyo7vei2OZM7pMI5ztxs/Q3DUU5RIQ/3gPQ/1E1IyQVsk3PrWDU
GOlWjH0W755pER6gJ4EucEbXI2Dhx15w+4N17JlFfAlz5xjj1E0iCQhWara4LQgPHK05T+W+YwX9
AWrJyhfy6enqDqjkHRuum7xxtKxwx1XgVdV+gs6MM0l+NmQCEQXMKuEnM7tPUw6klc7R6BtqebzO
KcBa9f4JGWLMLK8SoY2lkPc9Lz3nCC1/TmcSrqoeyjoMReUWPqCwPc7q6sD+wL8MAnMwEg9WjecU
hsUGJBlR6Fvyn/gzsK8cZwVpi5DcbZQgYYScgK0glQBkKsez54bct5UtxNqFPZDbNWxCwBclng21
pf1HebEML2dsAlSZv2UPWaHwGf3IiSwErkHynVCs/DfUWXdp5pPdCHQEDCvRoF8FZuIx10WflufS
bOfPRtUIJt8kj5n/pdsWUhfQBQd/q8Yz9LagWVReOah4Bu0O0UhTsxYT9iotWfC6mLJyK5BHRjWP
cILO3NAA6gQU2gRXIAnXRjQNBS4jks77OePHPeoR0rEagIoWzCh+3ce9sELMkeQEmL2NT7/J0I8H
52s2FaWrXI2pJeWt6X+DaFufl26naDlZo9TDlR86xx8/GRWghcjYGdYtfXVxxuaClY5vRRahktBA
1r5x6sDKdTFO/hsrTHlJjiTJUtPYGd6jD9wqUl+btYygfOq1RYIrqCrGkur+Xt0D06tz+vZxlC38
ZzWhorqvFprUsF2qEOrluYH3ILbqlgWzD31LWVGzcx8ZSQDE8B0XZpOABiaP0uODkwJrhztZUqMO
5Mr5Iq7zh+9ua+tpaW9gJE9I/VbIzlXcMyAplOMe2IxtFnnRwU4fqu9QfyoScVpPX224Pn8MMtdG
fLcvTfJDfdfwAdqTcYNpv+UDPG2jd9kSM4k+zPy/iVQBDSsipF1EnoRM+6G7eWgbjAM5bcmvNlBw
ZG7Et0F4DxSn7WI9yPHgp2hW9CTc/uiCbE0EhDer/rnZtHcwgYyUZ5tTVHyc9pQ70ksZp/bS7cew
VbcSSx0juV108rlNF1lS8pBiJjuiZgx5N0aKCh0JgkeDy6lhs1fRu9IazJhyO3aJVDnd47+zwdDL
NE2C72DXSCJHq/OE6w/j8ljAvbni+9o1T9wRuHpYj/z4obu0Gg/ZLGqvyFUjJUS+5Lrb1LExoc8X
X220Q8IJVsD3iT5Ayx7lZBxFtO0U+tmY6B8FT0Nku7uAeCmpTBYiRdmba6foRKyqLvI+IMrFVr6z
at0qsFG6vPwKzQrtrlSqLJ/BaWsw1U6R6TdQG555JLWrgkwmRYEDPouVwhZ0xzfBQTcANyF9QJBU
//0bxXYVZwM5+qIAD1JvVUu+lZQccKuXUeWbRGHQXUU8PRwBbM+j/YeZBPVN81honDhmP3A/l+I8
8KoEYiRgZHJxT9J+yVWQDWvDCFz3Qgi18wufNpq1D/KiABWN3YSgu7u+ZMQTwVJmVJWSIsNkYgPk
wIXC4kROcEFjPEUN4jPqiNSSqtcaWJoCvWBwxkPqRwmQsbCdNpuMr/kvMHXUQNXC2LaGRKZ3EZB6
rQj+H+lx9LwIxEh9U/N7hQLx8rkR9tdu8oFVVyMRLpSayvkIq2PMAvtK6afEDFLFdxfv7aWV3sO4
3+V0gzTKO/5lhnr6KiHBP+4046dcVjOOLY4jhRDSSx9bf2+FgMLohCKXTnCc6uMz0+76ONznCayY
sfTkXv5rcirs7YCzRiuA82DEJt5OVXqulIWwa7CwoBU4LuBI33pb+CJjE5/v1eAx+jsDdupwBY4f
xdeKmTtrW5k5+4cFlMMQ4IOEJHF+AILU8Om1HkAe3MaAHqfhQiIGSY902oO/kq49GLSB3crOukB7
vZ2OEDqgvuAZ+aZxzjapqi2ehHhu5bKwVzXIuohKKRCX95t6PAj9q4STQLb1rWaVaFOkgoGZ02PV
e7WwfUv0UMsRnD4WqZUhOS3AgJKqv6Y2sn1KzYiqYCv2t4OTjlv8fVTDpJFh6s24gPGmnm41KODv
2/fbUytrzf5tMV8HyZYl+gYyITkhDlmIxAsQGwR2cpMkYVGKdSEx3jtsy4Dj8L1WtOo369gnFsPa
dGgnQKjIuWdjOnzqb7EtsSKFCJ3u6Dl0DwhLWvZU8rCT6LkzA4n4DZ+Si/1XVqtCV8n+NZDDQmmg
eHCa5cgK356DcJkdHp2kkOF6vlKt0aku7Ota4RRNvvr9i+E+gHDoGqTA9qYWXPhSk7aqIghO49xE
x+3sXvEUYXHXZSiJTbiOHa79MbuhvoB4bO2mP5mdPPUGKTn/97RCxTM20ybn6JN8zb/3IN6qDytA
x43cC/TOCYh2SRJZ++IXFzmp4iqUQ6DrMpzqfmaNQjjtpLqHfZQWULXPVVoORIVzg7pkkg9QD4fs
ODmMkrRF6zBr7DHNFQYE4vA2ZT3QoITP8GvtzefcABIjdlYD3iOxDLQCbE7VK8VEJkCV3zCLsQPs
2qJN9yGkq05WjGMbfcOX3odaamxmPHmLlcvb12/PKTClreGy7L8Gf3y1m+qyQIx0951KhuPpurPy
AYzMF5kDairoHa0OCc06ylDJ+2635HBLLz3jQ2ad7oRuXnNKOVWOkN8tuG2KuTGb14yA9m7CWsJu
PrM9wrkolOy+/Ucxg/bwd3BOh2EhNpJIThG0RReHOthHF+KdVOnD9UmtwrlHpOw6QwJhy3P49wBK
IQcB9PNQkowzyUhVrdY9j6YsD9Qq74CuHJiytLvsmYIJBZjAwRSeIHVcP4PrsDVLnsqKT9CJQrXX
q3QSwKVXvc1qcIIFwFdyOpXrtCM2B/N+m+CmCicSDNB0s+97uEGssXxar7y93eX3D2r1vDdvTx4F
BYl3gMv3+Suu2rQTbXssOFJV0T3OmL1i8lWcWPL8UCWHIp7t0tllto8NcbygkbI6pzphwlZMpzkX
xzg7PB93o7FMvPzXSGlIxFQwbRNhliIX4HETnwqAIYnKnpCaCwvaILUr5OCnxMpYsQTimj5QQozf
dbozvvdF7DQCifkuyjpTCmNlC4XXalceGr/kUr7KtTyShOwarFsGnnN9lORqWhXH8VVudas5DDwx
oop2t0KLJc0ncuGq1o/v/0gIeSvF0iO6bT6e0viotridG6kmAgQ4zANLViB4zXxrdgLyzOq+bNJg
gPiBKeoRJznctdE8GcslkD9NoM2u7E7w2b+pPkqs5QGFTROEUMkDQciYhUtuWGHEr05p+XMWKCj3
Ll9wKk6rFTG5UB3sOMa3SpkzxsU6oa1rWXPSZNCpylhlQaPyIP/2COWahyipUJkUWd2SGCNf1rew
aw9FX/bkV3kfTw7T0wq1TEDtdS5j3wwyVKIk2GuxQ6UORodeTSM2Yeco8blpAVouBEKQluJU7B8u
lFZCvf1NVUfmpXPLhGZHoIHLyOno0w21HfbZPpS2+9mZv6V9N7f8YZJQOAlkdyrN1yWRqjb1dbe1
hP1dsPIDn9qoE/IV2z+42aT2gQhB8v8c5V+KPMivJrjXgduX+xCwYJclRM1v+M8MGR1n0y/ABqPC
zEU8VB6chYZuiRKUd9ZPuD98lOrwZsYiYw8978oAHZ0Er6QkdOodCAN1KYL3jIK6y7Nyfx88G00m
b173t6YTFYN0ivGipqu2uGSsV5G3IasgTJ8dK9b1MTK72jxDMAJrJWkWjcjc07ua7QqNbbDAoNoJ
M4IIsC9otvs6R2mJxpBhwHKH2tD2ORJaE1tG3oshantFVyWPBWpyLv5EUfDuOQSISGkcbkfPuYLj
KrJ0oYshjNm6jLetdfwz3IJP34wQfJQoFoo24xG+rq/DAWWhQ9UEcLysYluVjwDvMeYdkO4RHcXs
L/XgLecCM6IBh8rcKVxVy+z4AAHd4TwC2l991jyS2yj9nACdDPeg/hpDMLDAHt3Ey32wqsUvtnqu
CcwcnTPifHKdC0RBElWk1cQToEbSwaia5F6MnCJvS+4xCBlRzkngYieWcyIonhYHPRytdzX9uW9w
g83B11VVk9vJvMwMoO6QLCBZZEUva/nygO4GOzMyD3krvuwbzjJOD1jY2bBRRxbPuJjpvCaEl4N9
cJkoP1pV4PLNyxj0oYjskMhYGf86tgYqnQCCbNMKWdzDSCtX5UAf9s7405VTj1Fe3mZDkEJqc3Gv
hPh9SsQPo/fitD74LkJIM/20zqtFdW/qZ0/4DqdloNm9EFkccKaZqUQ5SNhJBxQ/PO7J5XSPRadx
4173NvT3yVakY68BAskftaFQGOcL4f6KxzXF5OTFdM6I8KOVpIepi2NTVsUvuZ1gC9jQkyQBUu85
DmbTZcy5oX6W5cwYt3t/i20QTrUaeYD8Yhczwt4q++OKteBwUB+BqAMf12640+Fx6UOyhPLw+VNu
tzFELPlKL9cC3lBlGlI9929wJjc95dS3MjA5QkJKlvARwO9uTzBIhRc5c5gMv4tFS8xwaM4Xz86S
1rOfeI1NwnFH8ZQjOX0ehyoIiAVU5zYsaYHL1+l1Ecns323nd8Kim2anIQzAMkGASV+FW8R4zxu/
KTN87xP0cu5W/ZrukxKZqrB9tNHLy4KqWNEbEp1g/pF+rL8F9I52ZCr44NTA1B76WHJyrDwF/OH3
6yRkNVcBF0bVlr1KfFhKF7akzfISU0DUsCabrK20Jz/iekHDVGhhwu/ZyGETA7A+NmXxBWmLkqew
ueknNVNa4Xgkg3cqmZnDGoajWk0WM5epegbXC52e5R7WxFFWTv+8C+kc4MsnOmbGaM7wbsh8hvFR
yr13g+BOKvAn1EsJoQpymXhAbwJ7OLHoEXiGdf2Kkinh7Mf2zLS+GArsRCFBPXKRxjaZlCVraUq6
KjnFo7sgN5SlMK6UlKeTIMk2KmeNYFsO1MHz90uGwd4a+gixtBipRnTUV8LBpOXqf3vNED7WbBYO
q40nXdJ0gXPzB6BVhw/PB0V0Fo53d4ZKjyoGw6VU7P0qwh8c5iXu38ehiEljicC+UzKndvhZZmrW
Ky7jy+nvqcz8YuJEYZnr1RkyqqwEDz6cu259Tz8XnnNustPMs93YzBzUK1ZrWw8gEX8pXAuQDwT1
Ij/+uRe13NrsukC4yCnrh0cVC3ZmQp5n3aXDXIRf6p2qwaD9spkXpBV06sGfhUrlhMmmImWiiRsm
g5lDAZCeDcRJFQyFeof2YHc7H/WXiFpAUR/3/jKrs4EuMpZNNvG+PVlE5itxeHh0gFc8MaSqzbSH
Kj42pG/W0KQYECJ7qQvQPveDA1K0yx+7soD7q88QgCE7P05h7bTRalx+j30MvGAqZ2MDtS0mpLHS
J/82y0qTmZPLwjlJBPoBY1KX5Wa2Xb4zKjb4zZdrouDPhoCgL+6cUBu6ouzSPpPzQr1dj6B1TeAl
l0uA44CkCG1cuunu4hbVD4ZkN6P5Kw03kt3DNMiEZoO45yneBn+a9RUZBEbTH5Se4InVVX/fQa7s
7CZ0rr7FLuTbLuaRqF5qMefvTKMXTywhH0Q8P3Xaz20N99hS0H11XR+8MaX9ljY7TUmuoegc0Usa
kTOR+47blwnP5W55Ip3ZFdcCnKzlV+vxon5UNK+t9QW67cQNg8imQzVzRIXugFaqlDN42PMTPZjy
l3bNucl+H+OBqmmZNdiRMDOPob1tF1rZZ7jQASA53J6tHUvq0rfiqCWJG3Q1oQYFehlgaWXsZe9R
pm8GGpncAfArxpfVT9HsOpf2TGd1B7mG+8+SzU0nro0dj8mjCNRgN7kCvB+gobD6hYA1/GNwP1rk
ZMOnopUBFC3GeydfWChpp4cZyBgQ/RDFoW/3Hrj448j34Fxl6YtHkJUmxNX4nsTBtlxwiu8OJWQT
ClDgrk/gebO9947XzQJE1GlpbVhfA+C0YD6/KTbZPTo5LsB8jvVF0v2sZdkJIL8xqfDbXQ==
`protect end_protected
